//================================================================================================
//    Date      Vers   Who  Changes
// -----------------------------------------------------------------------------------------------
// 17-Mar-2025  1.0.0  DWW  Initial creation
//================================================================================================
localparam VERSION_MAJOR = 1;
localparam VERSION_MINOR = 0;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 0;
localparam RTL_TYPE      = 31725;
localparam RTL_SUBTYPE   = 0;

localparam VERSION_DAY   = 17;
localparam VERSION_MONTH = 3;
localparam VERSION_YEAR  = 2025;
